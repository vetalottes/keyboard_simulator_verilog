`timescale 1ns / 1ps

module chars(
    input [5:0] char,
    input [2:0] rownum,
    output reg [7:0] pixels
    );
    
    initial pixels = 0;
    
    always@(*) begin
    case({char,rownum})
        9'b000000_000: pixels = 8'b01111100; // q
        9'b000000_001: pixels = 8'b10000010; 
        9'b000000_010: pixels = 8'b10000010; 
        9'b000000_011: pixels = 8'b10000010; 
        9'b000000_100: pixels = 8'b10001010; 
        9'b000000_101: pixels = 8'b01111100; 
        9'b000000_110: pixels = 8'b00000010;  
        9'b000000_111: pixels = 8'b00000000;         
                            
        9'b000001_000: pixels = 8'b10000010; // w
        9'b000001_001: pixels = 8'b10000010; 
        9'b000001_010: pixels = 8'b10000010; 
        9'b000001_011: pixels = 8'b10000010; 
        9'b000001_100: pixels = 8'b10000010; 
        9'b000001_101: pixels = 8'b01010100; 
        9'b000001_110: pixels = 8'b01101100;  
        9'b000001_111: pixels = 8'b00000000;  
        
        9'b000010_000: pixels = 8'b11111110; // e
        9'b000010_001: pixels = 8'b10000000; 
        9'b000010_010: pixels = 8'b10000000; 
        9'b000010_011: pixels = 8'b11111110; 
        9'b000010_100: pixels = 8'b10000000; 
        9'b000010_101: pixels = 8'b10000000; 
        9'b000010_110: pixels = 8'b11111110;  
        9'b000010_111: pixels = 8'b00000000;  
        
        9'b000011_000: pixels = 8'b11111100; // r
        9'b000011_001: pixels = 8'b10000010; 
        9'b000011_010: pixels = 8'b10000010; 
        9'b000011_011: pixels = 8'b11111100; 
        9'b000011_100: pixels = 8'b10001000; 
        9'b000011_101: pixels = 8'b10000100; 
        9'b000011_110: pixels = 8'b10000010;  
        9'b000011_111: pixels = 8'b00000000;  
        
        9'b000100_000: pixels = 8'b11111110; // t 
        9'b000100_001: pixels = 8'b10111010; 
        9'b000100_010: pixels = 8'b00111000; 
        9'b000100_011: pixels = 8'b00111000; 
        9'b000100_100: pixels = 8'b00111000; 
        9'b000100_101: pixels = 8'b00111000; 
        9'b000100_110: pixels = 8'b00111000;  
        9'b000100_111: pixels = 8'b00000000;  
        
        9'b000101_000: pixels = 8'b11000110; // y
        9'b000101_001: pixels = 8'b11000110; 
        9'b000101_010: pixels = 8'b11000110; 
        9'b000101_011: pixels = 8'b01101100; 
        9'b000101_100: pixels = 8'b00111000; 
        9'b000101_101: pixels = 8'b00111000; 
        9'b000101_110: pixels = 8'b00111000;  
        9'b000101_111: pixels = 8'b00000000;  
        
        9'b000110_000: pixels = 8'b10000010; // u 
        9'b000110_001: pixels = 8'b10000010; 
        9'b000110_010: pixels = 8'b10000010; 
        9'b000110_011: pixels = 8'b10000010; 
        9'b000110_100: pixels = 8'b10000010; 
        9'b000110_101: pixels = 8'b10000010; 
        9'b000110_110: pixels = 8'b01111100;  
        9'b000110_111: pixels = 8'b00000000;  
        
        9'b000111_000: pixels = 8'b11111110; // i 
        9'b000111_001: pixels = 8'b00111000; 
        9'b000111_010: pixels = 8'b00111000; 
        9'b000111_011: pixels = 8'b00111000; 
        9'b000111_100: pixels = 8'b00111000; 
        9'b000111_101: pixels = 8'b00111000; 
        9'b000111_110: pixels = 8'b11111110;  
        9'b000111_111: pixels = 8'b00000000;  
        
        9'b001000_000: pixels = 8'b01111100; // o 
        9'b001000_001: pixels = 8'b11000110; 
        9'b001000_010: pixels = 8'b11000110; 
        9'b001000_011: pixels = 8'b11000110; 
        9'b001000_100: pixels = 8'b11000110; 
        9'b001000_101: pixels = 8'b11000110; 
        9'b001000_110: pixels = 8'b01111100;  
        9'b001000_111: pixels = 8'b00000000;  
        
        9'b001001_000: pixels = 8'b11111100; // p 
        9'b001001_001: pixels = 8'b10000010; 
        9'b001001_010: pixels = 8'b10000010; 
        9'b001001_011: pixels = 8'b11111100; 
        9'b001001_100: pixels = 8'b10000000; 
        9'b001001_101: pixels = 8'b10000000; 
        9'b001001_110: pixels = 8'b10000000;  
        9'b001001_111: pixels = 8'b00000000;  
        
        9'b001010_000: pixels = 8'b00111100; // a 
        9'b001010_001: pixels = 8'b01000100; 
        9'b001010_010: pixels = 8'b10000010; 
        9'b001010_011: pixels = 8'b11111110; 
        9'b001010_100: pixels = 8'b10000010; 
        9'b001010_101: pixels = 8'b10000010; 
        9'b001010_110: pixels = 8'b10000010;  
        9'b001010_111: pixels = 8'b00000000;  
        
        9'b001011_000: pixels = 8'b01111000; // s 
        9'b001011_001: pixels = 8'b10000110; 
        9'b001011_010: pixels = 8'b10000000; 
        9'b001011_011: pixels = 8'b01111100; 
        9'b001011_100: pixels = 8'b00000010; 
        9'b001011_101: pixels = 8'b11000010; 
        9'b001011_110: pixels = 8'b00111100;  
        9'b001011_111: pixels = 8'b00000000;  
        
        9'b001100_000: pixels = 8'b11110000; // d 
        9'b001100_001: pixels = 8'b10001100; 
        9'b001100_010: pixels = 8'b10000010; 
        9'b001100_011: pixels = 8'b10000010; 
        9'b001100_100: pixels = 8'b10000010; 
        9'b001100_101: pixels = 8'b10001100; 
        9'b001100_110: pixels = 8'b11111000;  
        9'b001100_111: pixels = 8'b00000000;  
        
        9'b001101_000: pixels = 8'b11111110; // f 
        9'b001101_001: pixels = 8'b10000000; 
        9'b001101_010: pixels = 8'b10000000; 
        9'b001101_011: pixels = 8'b11111110; 
        9'b001101_100: pixels = 8'b10000000; 
        9'b001101_101: pixels = 8'b10000000; 
        9'b001101_110: pixels = 8'b10000000;  
        9'b001101_111: pixels = 8'b00000000;  
        
        9'b001110_000: pixels = 8'b00111000; // g 
        9'b001110_001: pixels = 8'b01000100; 
        9'b001110_010: pixels = 8'b10000000; 
        9'b001110_011: pixels = 8'b10000000; 
        9'b001110_100: pixels = 8'b10001100; 
        9'b001110_101: pixels = 8'b01000010; 
        9'b001110_110: pixels = 8'b00111100;  
        9'b001110_111: pixels = 8'b00000000;  
        
        9'b001111_000: pixels = 8'b11000110; // h 
        9'b001111_001: pixels = 8'b11000110; 
        9'b001111_010: pixels = 8'b11000110; 
        9'b001111_011: pixels = 8'b11111110; 
        9'b001111_100: pixels = 8'b11000110; 
        9'b001111_101: pixels = 8'b11000110; 
        9'b001111_110: pixels = 8'b11000110;  
        9'b001111_111: pixels = 8'b00000000;  
        
        9'b010000_000: pixels = 8'b00001110; // j 
        9'b010000_001: pixels = 8'b00000100; 
        9'b010000_010: pixels = 8'b00000100; 
        9'b010000_011: pixels = 8'b00000100; 
        9'b010000_100: pixels = 8'b00000100; 
        9'b010000_101: pixels = 8'b10000100; 
        9'b010000_110: pixels = 8'b11111000;  
        9'b010000_111: pixels = 8'b00000000;  
        
        9'b010001_000: pixels = 8'b10001000; // k 
        9'b010001_001: pixels = 8'b10010000; 
        9'b010001_010: pixels = 8'b10100000; 
        9'b010001_011: pixels = 8'b11000000; 
        9'b010001_100: pixels = 8'b10100000; 
        9'b010001_101: pixels = 8'b10010000; 
        9'b010001_110: pixels = 8'b10001000;  
        9'b010001_111: pixels = 8'b00000000;  
        
        9'b010010_000: pixels = 8'b01000000; // l 
        9'b010010_001: pixels = 8'b01000000; 
        9'b010010_010: pixels = 8'b01000000; 
        9'b010010_011: pixels = 8'b01000000; 
        9'b010010_100: pixels = 8'b01000000; 
        9'b010010_101: pixels = 8'b01000010; 
        9'b010010_110: pixels = 8'b01111110;  
        9'b010010_111: pixels = 8'b00000000;  
        
        9'b010011_000: pixels = 8'b11111110; // z 
        9'b010011_001: pixels = 8'b00000110; 
        9'b010011_010: pixels = 8'b00001000; 
        9'b010011_011: pixels = 8'b00010000; 
        9'b010011_100: pixels = 8'b00100000; 
        9'b010011_101: pixels = 8'b11000000; 
        9'b010011_110: pixels = 8'b11111110;  
        9'b010011_111: pixels = 8'b00000000;  
        
        9'b010100_000: pixels = 8'b10000010; // x 
        9'b010100_001: pixels = 8'b01000100; 
        9'b010100_010: pixels = 8'b00101000; 
        9'b010100_011: pixels = 8'b00010000; 
        9'b010100_100: pixels = 8'b00101000; 
        9'b010100_101: pixels = 8'b01000100; 
        9'b010100_110: pixels = 8'b10000010;  
        9'b010100_111: pixels = 8'b00000000;  
        
        9'b010101_000: pixels = 8'b00011110; // c 
        9'b010101_001: pixels = 8'b01100000; 
        9'b010101_010: pixels = 8'b11000000; 
        9'b010101_011: pixels = 8'b11000000; 
        9'b010101_100: pixels = 8'b11000000; 
        9'b010101_101: pixels = 8'b01100000; 
        9'b010101_110: pixels = 8'b00011110;  
        9'b010101_111: pixels = 8'b00000000;  
        
        9'b010110_000: pixels = 8'b10000010; // v 
        9'b010110_001: pixels = 8'b10000010; 
        9'b010110_010: pixels = 8'b01000100; 
        9'b010110_011: pixels = 8'b01000100; 
        9'b010110_100: pixels = 8'b00101000; 
        9'b010110_101: pixels = 8'b00101000; 
        9'b010110_110: pixels = 8'b00010000;  
        9'b010110_111: pixels = 8'b00000000;  
        
        9'b010111_000: pixels = 8'b11111100; // b 
        9'b010111_001: pixels = 8'b01100110; 
        9'b010111_010: pixels = 8'b01100110; 
        9'b010111_011: pixels = 8'b01111000; 
        9'b010111_100: pixels = 8'b01100110; 
        9'b010111_101: pixels = 8'b01100110; 
        9'b010111_110: pixels = 8'b11111100;  
        9'b010111_111: pixels = 8'b00000000;  
        
        9'b011000_000: pixels = 8'b10000010; // n 
        9'b011000_001: pixels = 8'b11000010; 
        9'b011000_010: pixels = 8'b10100010; 
        9'b011000_011: pixels = 8'b10010010; 
        9'b011000_100: pixels = 8'b10001010; 
        9'b011000_101: pixels = 8'b10000110; 
        9'b011000_110: pixels = 8'b10000010;  
        9'b011000_111: pixels = 8'b00000000;  
        
        9'b011001_000: pixels = 8'b10000010; // m 
        9'b011001_001: pixels = 8'b11000110; 
        9'b011001_010: pixels = 8'b10101010; 
        9'b011001_011: pixels = 8'b10010010; 
        9'b011001_100: pixels = 8'b10000010; 
        9'b011001_101: pixels = 8'b10000010; 
        9'b011001_110: pixels = 8'b10000010;  
        9'b011001_111: pixels = 8'b00000000; 
        
        9'b011010_000: pixels = 8'b11111110; // 0
        9'b011010_001: pixels = 8'b10000110; 
        9'b011010_010: pixels = 8'b10001010; 
        9'b011010_011: pixels = 8'b10010010; 
        9'b011010_100: pixels = 8'b10100010; 
        9'b011010_101: pixels = 8'b11000010; 
        9'b011010_110: pixels = 8'b11111110;  
        9'b011010_111: pixels = 8'b00000000;
        
        9'b011011_000: pixels = 8'b00000010; // 1
        9'b011011_001: pixels = 8'b00000110; 
        9'b011011_010: pixels = 8'b00001010; 
        9'b011011_011: pixels = 8'b00010010; 
        9'b011011_100: pixels = 8'b00000010; 
        9'b011011_101: pixels = 8'b00000010; 
        9'b011011_110: pixels = 8'b00000010;  
        9'b011011_111: pixels = 8'b00000000;
        
        9'b011100_000: pixels = 8'b11111110; // 2
        9'b011100_001: pixels = 8'b00000010; 
        9'b011100_010: pixels = 8'b00000010; 
        9'b011100_011: pixels = 8'b11111110; 
        9'b011100_100: pixels = 8'b10000000; 
        9'b011100_101: pixels = 8'b10000000; 
        9'b011100_110: pixels = 8'b11111110;  
        9'b011100_111: pixels = 8'b00000000;
        
        9'b011101_000: pixels = 8'b11111110; // 3
        9'b011101_001: pixels = 8'b00000010; 
        9'b011101_010: pixels = 8'b00000010; 
        9'b011101_011: pixels = 8'b11111110; 
        9'b011101_100: pixels = 8'b00000010; 
        9'b011101_101: pixels = 8'b00000010; 
        9'b011101_110: pixels = 8'b11111110;  
        9'b011101_111: pixels = 8'b00000000;
        
        9'b011110_000: pixels = 8'b10000010; // 4
        9'b011110_001: pixels = 8'b10000010; 
        9'b011110_010: pixels = 8'b10000010; 
        9'b011110_011: pixels = 8'b11111110; 
        9'b011110_100: pixels = 8'b00000010; 
        9'b011110_101: pixels = 8'b00000010; 
        9'b011110_110: pixels = 8'b00000010;  
        9'b011110_111: pixels = 8'b00000000;
        
        9'b011111_000: pixels = 8'b11111110; // 5
        9'b011111_001: pixels = 8'b10000000; 
        9'b011111_010: pixels = 8'b10000000; 
        9'b011111_011: pixels = 8'b11111110; 
        9'b011111_100: pixels = 8'b00000010; 
        9'b011111_101: pixels = 8'b00000010; 
        9'b011111_110: pixels = 8'b11111110;  
        9'b011111_111: pixels = 8'b00000000;
        
        9'b100000_000: pixels = 8'b11111110; // 6
        9'b100000_001: pixels = 8'b10000000; 
        9'b100000_010: pixels = 8'b10000000; 
        9'b100000_011: pixels = 8'b11111110; 
        9'b100000_100: pixels = 8'b10000010; 
        9'b100000_101: pixels = 8'b10000010; 
        9'b100000_110: pixels = 8'b11111110;  
        9'b100000_111: pixels = 8'b00000000;
        
        9'b100001_000: pixels = 8'b11111110; // 7
        9'b100001_001: pixels = 8'b00000100; 
        9'b100001_010: pixels = 8'b00001000; 
        9'b100001_011: pixels = 8'b00010000; 
        9'b100001_100: pixels = 8'b00100000; 
        9'b100001_101: pixels = 8'b01000000; 
        9'b100001_110: pixels = 8'b10000000;  
        9'b100001_111: pixels = 8'b00000000;
        
        9'b100010_000: pixels = 8'b11111110; // 8
        9'b100010_001: pixels = 8'b10000010; 
        9'b100010_010: pixels = 8'b10000010; 
        9'b100010_011: pixels = 8'b11111110; 
        9'b100010_100: pixels = 8'b10000010; 
        9'b100010_101: pixels = 8'b10000010; 
        9'b100010_110: pixels = 8'b11111110;  
        9'b100010_111: pixels = 8'b00000000;
        
        9'b100011_000: pixels = 8'b11111110; // 9
        9'b100011_001: pixels = 8'b10000010; 
        9'b100011_010: pixels = 8'b10000010; 
        9'b100011_011: pixels = 8'b11111110; 
        9'b100011_100: pixels = 8'b00000010; 
        9'b100011_101: pixels = 8'b00000010; 
        9'b100011_110: pixels = 8'b11111110;  
        9'b100011_111: pixels = 8'b00000000;
        
        9'b100100_000: pixels = 8'b00000000; // ,
        9'b100100_001: pixels = 8'b00000000; 
        9'b100100_010: pixels = 8'b00000000; 
        9'b100100_011: pixels = 8'b00000000; 
        9'b100100_100: pixels = 8'b01100000; 
        9'b100100_101: pixels = 8'b00010000; 
        9'b100100_110: pixels = 8'b00100000;  
        9'b100100_111: pixels = 8'b00000000;
        
        9'b100101_000: pixels = 8'b00000000; // .
        9'b100101_001: pixels = 8'b00000000; 
        9'b100101_010: pixels = 8'b00000000; 
        9'b100101_011: pixels = 8'b00000000; 
        9'b100101_100: pixels = 8'b00000000; 
        9'b100101_101: pixels = 8'b00111000; 
        9'b100101_110: pixels = 8'b00111000;  
        9'b100101_111: pixels = 8'b00000000;
        
        9'b100110_000: pixels = 8'b00000010; // /
        9'b100110_001: pixels = 8'b00000100; 
        9'b100110_010: pixels = 8'b00001000; 
        9'b100110_011: pixels = 8'b00010000; 
        9'b100110_100: pixels = 8'b00100000; 
        9'b100110_101: pixels = 8'b01000000; 
        9'b100110_110: pixels = 8'b10000000;  
        9'b100110_111: pixels = 8'b00000000;
        
        9'b100111_000: pixels = 8'b00000000; // ;
        9'b100111_001: pixels = 8'b00110000; 
        9'b100111_010: pixels = 8'b00110000; 
        9'b100111_011: pixels = 8'b00000000; 
        9'b100111_100: pixels = 8'b00110000; 
        9'b100111_101: pixels = 8'b00001000; 
        9'b100111_110: pixels = 8'b00010000;  
        9'b100111_111: pixels = 8'b00000000;
        
        9'b101000_000: pixels = 8'b00001000; // '
        9'b101000_001: pixels = 8'b00001000; 
        9'b101000_010: pixels = 8'b00001000; 
        9'b101000_011: pixels = 8'b00000000; 
        9'b101000_100: pixels = 8'b00000000; 
        9'b101000_101: pixels = 8'b00000000; 
        9'b101000_110: pixels = 8'b00000000;  
        9'b101000_111: pixels = 8'b00000000;
        
        9'b101001_000: pixels = 8'b00000000; // -
        9'b101001_001: pixels = 8'b00000000; 
        9'b101001_010: pixels = 8'b00000000; 
        9'b101001_011: pixels = 8'b11111110; 
        9'b101001_100: pixels = 8'b00000000; 
        9'b101001_101: pixels = 8'b00000000; 
        9'b101001_110: pixels = 8'b00000000;  
        9'b101001_111: pixels = 8'b00000000;
        
        9'b101010_000: pixels = 8'b00000000; // =
        9'b101010_001: pixels = 8'b00000000; 
        9'b101010_010: pixels = 8'b11111110; 
        9'b101010_011: pixels = 8'b00000000; 
        9'b101010_100: pixels = 8'b11111110; 
        9'b101010_101: pixels = 8'b00000000; 
        9'b101010_110: pixels = 8'b00000000;  
        9'b101010_111: pixels = 8'b00000000;
        
        9'b101011_000: pixels = 8'b11110000; // [
        9'b101011_001: pixels = 8'b10000000; 
        9'b101011_010: pixels = 8'b10000000; 
        9'b101011_011: pixels = 8'b10000000; 
        9'b101011_100: pixels = 8'b10000000; 
        9'b101011_101: pixels = 8'b10000000; 
        9'b101011_110: pixels = 8'b11110000;  
        9'b101011_111: pixels = 8'b00000000;
        
        9'b101100_000: pixels = 8'b00011110; // ]
        9'b101100_001: pixels = 8'b00000010; 
        9'b101100_010: pixels = 8'b00000010; 
        9'b101100_011: pixels = 8'b00000010; 
        9'b101100_100: pixels = 8'b00000010; 
        9'b101100_101: pixels = 8'b00000010; 
        9'b101100_110: pixels = 8'b00011110;  
        9'b101100_111: pixels = 8'b00000000;
        
        9'b101101_000: pixels = 8'b10000000; // \
        9'b101101_001: pixels = 8'b01000000; 
        9'b101101_010: pixels = 8'b00100000; 
        9'b101101_011: pixels = 8'b00010000; 
        9'b101101_100: pixels = 8'b00001000; 
        9'b101101_101: pixels = 8'b00000100; 
        9'b101101_110: pixels = 8'b00000010;  
        9'b101101_111: pixels = 8'b00000000; 
        
        9'b111111_000: pixels = 8'b00000000; // null
        9'b111111_001: pixels = 8'b00000000; 
        9'b111111_010: pixels = 8'b00000000;     
        9'b111111_011: pixels = 8'b00000000;    
        9'b111111_100: pixels = 8'b00000000;     
        9'b111111_101: pixels = 8'b00000000;    
        9'b111111_110: pixels = 8'b00000000;    
        9'b111111_111: pixels = 8'b00000000; 
        default: pixels = 8'b00000000;
   endcase
   end
endmodule
